package interfaces;
    `include "interfaces.svh"
endpackage

package structs_and_typedefs;
    `include "structs_and_typedefs.svh"
endpackage

package parameters;
    `include "parameters.svh"
endpackage

